-------------------------------------------------------------------------------
-- Module     : t_traffic_light_phase_cnt
-------------------------------------------------------------------------------
-- Author     : <haf@fh-augsburg.de>
-- Company    : University of Applied Sciences Augsburg
-- Copyright (c) 2011   <haf@fh-augsburg.de>
-------------------------------------------------------------------------------
-- Description: Testbench for design "traffic_light_phase_cnt"
-------------------------------------------------------------------------------
-- Revisions  : see end of file
-------------------------------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY t_traffic_light_phase_cnt IS
END t_traffic_light_phase_cnt;

ARCHITECTURE tbench OF t_traffic_light_phase_cnt IS

  COMPONENT traffic_light IS
    PORT (
      clk             : IN  std_ulogic;
      rst_n           : IN  std_ulogic;
      en_pi           : IN  std_ulogic;
      end_of_phase_pi : IN  std_ulogic;
      ld_cnt_po       : OUT std_ulogic;
      phase_select_o  : OUT std_ulogic_vector(1 DOWNTO 0);
      ns_red_o        : OUT std_ulogic;
      ns_yellow_o     : OUT std_ulogic;
      ns_green_o      : OUT std_ulogic;
      ew_red_o        : OUT std_ulogic;
      ew_yellow_o     : OUT std_ulogic;
      ew_green_o      : OUT std_ulogic);
  END COMPONENT traffic_light;
  
  -- definition of a clock period
  CONSTANT period : time    := 20 ns;
  -- switch for clock generator
  SIGNAL clken_p  : boolean := true;


  -- component ports
  SIGNAL clk_i           : std_ulogic;
  SIGNAL rst_ni          : std_ulogic;
  SIGNAL red_phase_value : std_ulogic_vector(3 DOWNTO 0);
  SIGNAL ry_phase_value  : std_ulogic_vector(3 DOWNTO 0);
  SIGNAL g_phase_value   : std_ulogic_vector(3 DOWNTO 0);
  SIGNAL y_phase_value   : std_ulogic_vector(3 DOWNTO 0);
  SIGNAL count_o         : std_ulogic_vector(3 DOWNTO 0);
  SIGNAL ns_red_o        : std_ulogic;
  SIGNAL ns_yellow_o     : std_ulogic;
  SIGNAL ns_green_o      : std_ulogic;
  SIGNAL ew_red_o        : std_ulogic;
  SIGNAL ew_yellow_o     : std_ulogic;
  SIGNAL ew_green_o      : std_ulogic;
  
  SIGNAL scaled_period : std_ulogic;

BEGIN  -- tbench

  -- component instantiation
  DUT : ENTITY work.traffic_light_phase_cnt(structure)
    PORT MAP (
      clk_i           => clk_i,
      rst_ni          => rst_ni,
      en_pi           => scaled_period,
      red_phase_value => red_phase_value,
      ry_phase_value  => ry_phase_value,
      g_phase_value   => g_phase_value,
      y_phase_value   => y_phase_value,
      count_o         => count_o,
      ns_red_o        => ns_red_o,
      ns_yellow_o     => ns_yellow_o,
      ns_green_o      => ns_green_o,
      ew_red_o        => ew_red_o,
      ew_yellow_o     => ew_yellow_o,
      ew_green_o      => ew_green_o);
 
  -- clock generation
  clock_proc : PROCESS
  BEGIN
    WHILE clken_p LOOP
      clk_i <= '0'; WAIT FOR period/2;
      clk_i <= '1'; WAIT FOR period/2;
    END LOOP;
    WAIT;
  END PROCESS;

  -- initial reset, always necessary at the beginning of a simulation
  reset : rst_ni <= '0', '1' AFTER period;

  ---------------------------------------------------------------------
  -- prescaler, generates an enable signal
  -- in dependence of clock period and generic parameter m
  clock_divider : ENTITY work.cntdnmodm(rtl)
    GENERIC MAP (
      n => 3,
      m => 4)
    PORT MAP (
      clk_i   => clk_i,
      rst_ni  => rst_ni,
      en_pi   => '1',                   -- permanently enabled
      count_o => OPEN,                  -- open, because not needed
      tc_o    => scaled_period);
  ---------------------------------------------------------------------

  stimuli_p : PROCESS

  BEGIN

    WAIT UNTIL rst_ni = '1';            -- wait until asynchronous reset ...
                                        -- ... is deactivated

    ---------------------------------------------------------------------------
    red_phase_value <= "0101";          -- set phase values
    ry_phase_value  <= "0000";
    g_phase_value   <= X"3";  
    y_phase_value   <= X"0";  

    WAIT FOR 900 ns;                    -- wait for at least a full cycle
    ---------------------------------------------------------------------------

    -- Follow the comments below to continue verification
    ---------------------------------------------------------------------------
              -- change red phase value
    
    
              -- change green phase value
    
    
              -- wait for at least a full cycle
    ---------------------------------------------------------------------------
    
    

    clken_p <= false;                   -- switch clock generator off

    WAIT;
  END PROCESS;

END tbench;

-------------------------------------------------------------------------------
-- Revisions:
-- ----------
-- $Id:$
-------------------------------------------------------------------------------
