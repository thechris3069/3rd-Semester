-------------------------------------------------------------------------------
-- Module     : t_traffic_light
-------------------------------------------------------------------------------
-- Author     : <haf@fh-augsburg.de>
-- Company    : University of Applied Sciences Augsburg
-- Copyright (c) 2011   <haf@fh-augsburg.de>
-------------------------------------------------------------------------------
-- Description: Testbench for design "traffic_light"
-------------------------------------------------------------------------------
-- Revisions  : see end of file
-------------------------------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY t_traffic_light IS
END t_traffic_light;

ARCHITECTURE tbench OF t_traffic_light IS
  COMPONENT traffic_light IS
    PORT (
      clk              : IN  std_ulogic;
      rst_n            : IN  std_ulogic;
      next_phase_en_pi : IN  std_ulogic;
      red_o            : OUT std_ulogic;
      yellow_o         : OUT std_ulogic;
      green_o          : OUT std_ulogic);
  END COMPONENT traffic_light;
  
  -- definition of a clock period
  CONSTANT period : time    := 20 ns;
  -- switch for clock generator
  SIGNAL clken_p  : boolean := true;


  -- component ports
  SIGNAL clk_i           : std_ulogic;
  SIGNAL rst_ni          : std_ulogic;

  SIGNAL red_o            : std_ulogic;
  SIGNAL yellow_o         : std_ulogic;
  SIGNAL green_o          : std_ulogic;
   
  SIGNAL scaled_period : std_ulogic;

BEGIN  -- tbench
  
  -- component instantiation
  DUT : ENTITY work.traffic_light
    PORT MAP (
      clk              => clk_i,
      rst_n            => rst_ni,
      next_phase_en_pi => scaled_period,
      red_o            => red_o,
      yellow_o         => yellow_o,
      green_o          => green_o);
 
  -- clock generation
  clock_proc : PROCESS
  BEGIN
    WHILE clken_p LOOP
      clk_i <= '0'; WAIT FOR period/2;
      clk_i <= '1'; WAIT FOR period/2;
    END LOOP;
    WAIT;
  END PROCESS;

  -- initial reset, always necessary at the beginning of a simulation
  reset : rst_ni <= '0', '1' AFTER period;

  ---------------------------------------------------------------------
  -- prescaler, generates an enable signal
  -- in dependence of clock period and generic parameter m
  clock_divider : ENTITY work.cntdnmodm(rtl)
    GENERIC MAP (
      n => 3,
      m => 4)
    PORT MAP (
      clk_i   => clk_i,
      rst_ni  => rst_ni,
      en_pi   => '1',                   -- permanently enabled
      count_o => OPEN,                  -- open, because not needed
      tc_o    => scaled_period);
  ---------------------------------------------------------------------

  stimuli_p : PROCESS

  BEGIN

    WAIT UNTIL rst_ni = '1';            -- wait until asynchronous reset ...
                                        -- ... is deactivated

    ---------------------------------------------------------------------------
    
    WAIT FOR 800 ns;                    -- for at least a full cycle
    ---------------------------------------------------------------------------

    

    clken_p <= false;                   -- switch clock generator off

    WAIT;
  END PROCESS;

END tbench;

-------------------------------------------------------------------------------
-- Revisions:
-- ----------
-- $Id:$
-------------------------------------------------------------------------------
