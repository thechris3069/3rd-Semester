-------------------------------------------------------------------------------
-- Module     : t_add4
-------------------------------------------------------------------------------
-- Author     :   <haf@fh-augsburg.de>
-- Company    : University of Applied Sciences Augsburg
-- Copyright (c) 2011   <haf@fh-augsburg.de>
-------------------------------------------------------------------------------
-- Description: Testbench for design "add4"
-------------------------------------------------------------------------------
-- Revisions  : see end of file
-------------------------------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-------------------------------------------------------------------------------

ENTITY t_add4 IS
END t_add4;

-------------------------------------------------------------------------------

ARCHITECTURE tbench OF t_add4 IS

  COMPONENT add4
    PORT (
      a_i   : IN  std_ulogic_vector(3 DOWNTO 0);
      b_i   : IN  std_ulogic_vector(3 DOWNTO 0);
      ci_i  : IN  std_ulogic;
      sum_o : OUT std_ulogic_vector(3 DOWNTO 0);
      co_o  : OUT std_ulogic);
  END COMPONENT;

  -- definition of a clock period
  CONSTANT period : time := 10 ns;

  -- component ports
  SIGNAL a_i   : std_ulogic_vector(3 DOWNTO 0);
  SIGNAL b_i   : std_ulogic_vector(3 DOWNTO 0);
  SIGNAL ci_i  : std_ulogic;
  SIGNAL sum_o : std_ulogic_vector(3 DOWNTO 0);
  SIGNAL co_o  : std_ulogic;

BEGIN  -- tbench

  -- component instantiation
  DUT : ENTITY work.add4(structure)
    PORT MAP (
      a_i   => a_i,
      b_i   => b_i,
      ci_i  => ci_i,
      sum_o => sum_o,
      co_o  => co_o);

  stimuli_p : PROCESS

    -- purpose: apply stimuli to input signals of module under test
    PROCEDURE apply_stimuli (
      CONSTANT ci_stim        : IN std_ulogic;
      CONSTANT b_stim, a_stim : IN std_ulogic_vector) IS
    BEGIN  -- apply_stimuli
      a_i  <= a_stim;
      b_i  <= b_stim;
      ci_i <= ci_stim;
      WAIT FOR period;
    END PROCEDURE apply_stimuli;
  
  BEGIN
    a_i  <= X"0";            -- set a value to input a_i as hexadecimal value
    b_i  <= B"0000";         -- set a value to input b_i as binary vector value
    ci_i <= '0';             -- set a value to input ci_i as a 1-bit value
    WAIT FOR period;         -- values are assigned here

                             -- prefix B is the default, hence not necessary to write
    a_i <= "1111";           -- change value of a_i as binary vector value
    WAIT FOR period;

    a_i <= X"0";             -- change value of a_i
    b_i <= X"F";             -- change value of b_i
    WAIT FOR period;

    -- add your stimuli here ...

  apply_stimuli('1', X"1", X"0");
  apply_stimuli('1', X"1", X"1");
  apply_stimuli('1', X"1", X"2");
  apply_stimuli('1', X"0", X"2");
  apply_stimuli('1', X"0", X"F");
  
  apply_stimuli('1', X"5", X"E");
  
  apply_stimuli('0', X"5", X"E");
  
	
    -- alternatively, a local procedure can be used to assign input values:
	-----------------------------------------------------------------------
--                  ci_i, b_i,    a_i
    --apply_stimuli('0', B"0000", X"0");
    --apply_stimuli('0', B"1111", X"0");
    --apply_stimuli('0', X"F",    X"0");

    -- add your stimuli here ...

    
    WAIT;
  END PROCESS;

END tbench;

-------------------------------------------------------------------------------
-- Revisions:
-- ----------
-- $Id:$
-------------------------------------------------------------------------------
